module Main(input i_Clk);
endmodule
